module not_gate_primitive (
       input wire a,
       output wire y
   );
       not (y, a);
endmodule