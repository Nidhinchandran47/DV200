module not_gate_assign (
       input wire a,
       output wire y
   );
       assign y = ~a;
endmodule