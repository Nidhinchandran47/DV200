module and_gate_primitive (
    input wire a,
    input wire b,
    output wire y
);
    and (y, a, b);
endmodule
